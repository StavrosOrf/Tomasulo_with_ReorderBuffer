library IEEE;
use IEEE.STD_LOGIC_1164.all;

package my_Package_VectorV is

type Array_of_RegV is array(0 to 31) of std_logic_vector (31 downto 0);


end my_Package_VectorV;

